module NOT_gate_level(output Y, input A);
    not (Y, A);
endmodule